Linear Circuit

R1 1 2 500
C1 3 0 10n
L1 2 3 10m
Vb 1 0 AC 1
.AC DEC 100 1 100meg
.End
